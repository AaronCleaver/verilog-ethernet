/*

Copyright (c) 2016-2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * Generic ODDR module
 */
module oddr #
(
    // target ("SIM", "GENERIC", "XILINX", "ALTERA")
    parameter TARGET = "GENERIC",
    // IODDR style ("IODDR", "IODDR2")
    // Use IODDR for Virtex-4, Virtex-5, Virtex-6, 7 Series, Ultrascale
    // Use IODDR2 for Spartan-6
    parameter IODDR_STYLE = "IODDR2",
    // Width of register in bits
    parameter WIDTH = 1
)
(
    input  wire             clk,

    input  wire [WIDTH-1:0] d1,
    input  wire [WIDTH-1:0] d2,

    output wire [WIDTH-1:0] q
);

/*

Provides a consistent output DDR flip flop across multiple FPGA families
              _____       _____       _____       _____
    clk  ____/     \_____/     \_____/     \_____/     \_____
         _ ___________ ___________ ___________ ___________ __
    d1   _X____D0_____X____D2_____X____D4_____X____D6_____X__
         _ ___________ ___________ ___________ ___________ __
    d2   _X____D1_____X____D3_____X____D5_____X____D7_____X__
         _____ _____ _____ _____ _____ _____ _____ _____ ____
    d    _____X_D0__X_D1__X_D2__X_D3__X_D4__X_D5__X_D6__X_D7_

*/

genvar n;

generate

if (TARGET == "XILINX") begin
    for (n = 0; n < WIDTH; n = n + 1) begin : oddr
        if (IODDR_STYLE == "IODDR") begin
            ODDR #(
                .DDR_CLK_EDGE("SAME_EDGE"),
                .SRTYPE("ASYNC")
            )
            oddr_inst (
                .Q(q[n]),
                .C(clk),
                .CE(1'b1),
                .D1(d1[n]),
                .D2(d2[n]),
                .R(1'b0),
                .S(1'b0)
            );
        end else if (IODDR_STYLE == "IODDR2") begin
            ODDR2 #(
                .DDR_ALIGNMENT("C0"),
                .SRTYPE("ASYNC")
            )
            oddr_inst (
                .Q(q[n]),
                .C0(clk),
                .C1(~clk),
                .CE(1'b1),
                .D0(d1[n]),
                .D1(d2[n]),
                .R(1'b0),
                .S(1'b0)
            );
        end
    end
end else if (TARGET == "ALTERA") begin
    altddio_out #(
        .WIDTH(WIDTH),
        .POWER_UP_HIGH("OFF"),
        .OE_REG("UNUSED")
    )
    altddio_out_inst (
        .aset(1'b0),
        .datain_h(d1),
        .datain_l(d2),
        .outclocken(1'b1),
        .outclock(clk),
        .aclr(1'b0),
        .dataout(q)
    );
end else if (TARGET == "ALTERA_MAX10") begin
    altera_gpio_lite #(
      .PIN_TYPE                                 ("output"),
      .SIZE                                     (WIDTH),
      .REGISTER_MODE                            ("ddr"),
      .BUFFER_TYPE                              ("single-ended"),
      .ASYNC_MODE                               ("none"),
      .SYNC_MODE                                ("none"),
      .BUS_HOLD                                 ("false"),
      .OPEN_DRAIN_OUTPUT                        ("false"),
      .ENABLE_OE_PORT                           ("false"),
      .ENABLE_NSLEEP_PORT                       ("false"),
      .ENABLE_CLOCK_ENA_PORT                    ("false"),
      .SET_REGISTER_OUTPUTS_HIGH                ("false"),
      .INVERT_OUTPUT                            ("false"),
      .INVERT_INPUT_CLOCK                       ("false"),
      .USE_ONE_REG_TO_DRIVE_OE                  ("false"),
      .USE_DDIO_REG_TO_DRIVE_OE                 ("false"),
      .USE_ADVANCED_DDR_FEATURES                ("false"),
      .USE_ADVANCED_DDR_FEATURES_FOR_INPUT_ONLY ("false"),
      .ENABLE_OE_HALF_CYCLE_DELAY               ("true"),
      .INVERT_CLKDIV_INPUT_CLOCK                ("false"),
      .ENABLE_PHASE_INVERT_CTRL_PORT            ("false"),
      .ENABLE_HR_CLOCK                          ("false"),
      .INVERT_OUTPUT_CLOCK                      ("false"),
      .INVERT_OE_INCLOCK                        ("false"),
      .ENABLE_PHASE_DETECTOR_FOR_CK             ("false")
    ) max10_oddr_inst (
      .outclock        (clk), // outclock.export
      .din             ({d2,d1}),      //      din.export
      .pad_out         (q),  //  pad_out.export
      .outclocken      (1'b1),     // (terminated)
      .inclock         (1'b0),     // (terminated)
      .inclocken       (1'b0),     // (terminated)
      .fr_clock        (),         // (terminated)
      .hr_clock        (),         // (terminated)
      .invert_hr_clock (1'b0),     // (terminated)
      .phy_mem_clock   (1'b0),     // (terminated)
      .mimic_clock     (),         // (terminated)
      .dout            (),         // (terminated)
      .pad_io          (),         // (terminated)
      .pad_io_b        (),         // (terminated)
      .pad_in          ({WIDTH{1'b0}}),     // (terminated)
      .pad_in_b        ({WIDTH{1'b0}}),     // (terminated)
      .pad_out_b       (),         // (terminated)
      .aset            (1'b0),     // (terminated)
      .aclr            (1'b0),     // (terminated)
      .sclr            (1'b0),     // (terminated)
      .nsleep          ({WIDTH{1'b0}}),     // (terminated)
      .oe              ({WIDTH{1'b0}})      // (terminated)
    );
end else begin
    reg [WIDTH-1:0] d_reg_1 = {WIDTH{1'b0}};
    reg [WIDTH-1:0] d_reg_2 = {WIDTH{1'b0}};

    reg [WIDTH-1:0] q_reg = {WIDTH{1'b0}};

    always @(posedge clk) begin
        d_reg_1 <= d1;
        d_reg_2 <= d2;
    end

    always @(posedge clk) begin
        q_reg <= d1;
    end

    always @(negedge clk) begin
        q_reg <= d_reg_2;
    end

    assign q = q_reg;
end

endgenerate

endmodule
